module IM(input [15:0] addr,output [31:0] out_ins);
    reg [31:0] memory [0:255];
    reg [31:0] out_ins;
    integer i;
    initial begin
        for(i=0;i<=255;i=i+1) begin
            memory[i]=0;
        end
        memory[0]=32'b00000100000100000000000000000000; //reg0=reg2+reg1=3
        memory[1]=32'b00000000000100100000000000000001; //reg4=reg0-reg1=2
        memory[2]=32'b00011000001100000000000000010100; //reg0=reg12&reg30=0
        memory[3]=32'b10000000000000000000000010000000; //reg0+=8=8
        memory[4]=32'b10000000000000000000000001000011; //reg0/=4=2
        memory[5]=32'b10000010000000000000000000101011; //reg1=2
        memory[6]=32'b10000010000000000000000000001100; //DM[0]=reg1=2
        memory[7]=32'b01000010011100000000000000001000; //DM[reg7(7)]=reg1=2
        memory[8]=32'b10001100000000000000001100001010; //reg6=DM[48]=48
        memory[9]=32'b10000000000000000000000000101011; //reg0=2
        memory[10]=32'b01000000000100000000000000100001; //reg0==reg1?->PC+=2(=12)(triggered)
        //memory[10]=32'b01000000000100000000000011000000; //reg0==reg1?->PC=12(triggered)
        memory[11]=32'b01000000000100000000000000100001; //reg0==reg1?->PC+=2(skipped)
        memory[12]=32'b00000100000100000000000000000000; //reg2+reg1->reg0=4
        memory[13]=32'b01000000000100000000000000100010; //reg0==reg1?->PC=DM[2]=2(untriggered)
        //memory[14]=32'b01000100000100000000000001000010; //reg2==reg1?->PC=DM[4]=4(triggered)
        //memory[14]=32'b11000000000000000000000001000000; //jmp 4
        //memory[14]=32'b10000000000000000000000000001101; //jmp (reg0=4)
        memory[14]=32'b10000100000000000000000000101110; //jmp (reg3+2=4)
        memory[15]=32'b11000000000000000000000001010011; //PC+=DM[5](=9)(invalid)
    end
    always@(*)begin
        out_ins=memory[addr];
    end
endmodule